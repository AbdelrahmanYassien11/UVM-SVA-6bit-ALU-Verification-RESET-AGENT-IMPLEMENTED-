package rst_uvm_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"
/************************************
***********Sequence Items********
************************************/
`include "rst_sequence_item.sv"

/************************************
**********ALU Agent Components*******
************************************/
`include "rst_driver.sv"
`include "rst_monitor.sv"
`include "rst_sequencer.sv"

/************************************
*************Agents Configs**********
************************************/
`include "rst_agnt_cfg.sv"

/************************************
********Environment Components******
************************************/
`include "rst_agent.sv"

endpackage : rst_uvm_pkg